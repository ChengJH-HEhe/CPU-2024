`include "const.v"

// 8:2
module Bpredictor (
  input wire                 clk_in,			// system clock signal
  input wire                 rst_in,			// reset signal
  input wire					rdy_in,			// ready signal, pause cpu when low

  // insfetcher ask for prediction
  input wire [31 : 0] input_ins,
  input wire [31 : 0] input_pc,
  output wire predict_jump,
  output wire [31 : 0] predict_pc,

  // ROB update predictor
  input wire ROB_valid,
  input wire [31 : 0] ins_pc,
  input wire success
);
  localparam RISC_B = 7'b1100011;
  reg [1:0] state[127:0];

assign predict_jump = input_ins[6:0] == RISC_B? state[input_pc[8:2]][1] : 1'b0;
assign predict_pc = predict_jump? input_pc + {{20{input_ins[31]}},input_ins[7], input_ins[30:25], input_ins[11:8], 1'b0} : input_pc + 4;

integer i;
always @(posedge clk_in) begin
  if(rst_in) begin
    for(i = 0; i < 128; i = i + 1) begin
      state[i] <= 2'b00;
    end
  end else begin
    if(ROB_valid) 
      begin
        if(success) begin
          if(state[ins_pc[8:2]] != 2'b11)
            state[ins_pc[8:2]] <=   state[ins_pc[8:2]] + 1;
        end else begin
          if(state[ins_pc[8:2]] != 2'b00)
            state[ins_pc[8:2]] <=   state[ins_pc[8:2]] - 1;
        end
    end
  end
end
endmodule